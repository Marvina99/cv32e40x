module scoreboard import cv32e40x_pkg::*; 
#(
    //parameters
) 
(
    input scoreboard_entries_t scoreboard_entries__id_i,
    input scoreboard_entries_t scoreboard_entries__ex_i,
    input scoreboard_entries_t scoreboard_entries__lsu_i,
    input scoreboard_entries_t scoreboard_entries__wb_i
);
    
endmodule